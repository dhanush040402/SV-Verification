interface intr;
  logic a;
  logic b;
  logic sum;
  logic carry;
endinterface
